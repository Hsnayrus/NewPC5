module dffe(p]